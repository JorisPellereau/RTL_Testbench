//                              -*- Mode: Verilog -*-
// Filename        : pkg_tb.sv
// Description     : Testbench Package
// Author          : Linux-JP
// Created On      : Thu Sep 21 18:36:48 2023
// Last Modified By: Linux-JP
// Last Modified On: Thu Sep 21 18:36:48 2023
// Update Count    : 0
// Status          : Unknown, Use with caution!

package pkg_tb;

`include "tb_utils_class.sv"
`include "tb_set_injector_class.sv"
`include "tb_wait_event_class.sv"
`include "tb_check_level_class.sv"
`include "tb_modelsim_cmd_class.sv"
`include "tb_uart_class.sv"
`include "tb_data_collector_class.sv"
`include "tb_data_checker_class.sv"
`include "tb_master_axi4lite_class.sv"
`include "tb_i2c_slave_class.sv"

// TB Modules Custom Class contains previous class, so it is declare in last position
`include "tb_modules_custom_class.sv"

   
endpackage // pkg_tb
